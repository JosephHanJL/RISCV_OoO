/////////////////////////////////////////////////////////////////////////
//                                                                     //
//   Modulename :  vtuber_test.sv                                      //
//                                                                     //
//  Description :  Visual Debugger for project 4                       //
//                 Outputs only IF part                                //
//                                                                     //
/////////////////////////////////////////////////////////////////////////


`include "verilog/sys_defs.svh"

extern void initcurses(int,int,int,int,int,int,int,int,int,int);
extern void flushpipe();
extern void waitforresponse();
extern void initmem();
extern int get_instr_at_pc(int);
extern int not_valid_pc(int);

module testbench;
    string program_memory_file;

    // Registers and wires used in the testbench
    logic        clock;
    logic        reset;
    logic [31:0] clock_count;
    logic [31:0] instr_count;
    int          wb_fileno;
    logic [63:0] debug_counter; // counter used for when pipeline infinite loops, forces termination

    logic [1:0]       proc2mem_command;
    logic [`XLEN-1:0] proc2mem_addr;
    logic [63:0]      proc2mem_data;
    logic [3:0]       mem2proc_response;
    logic [63:0]      mem2proc_data;
    logic [3:0]       mem2proc_tag;
`ifndef CACHE_MODE
    MEM_SIZE          proc2mem_size;
`endif

    logic [3:0]            pipeline_completed_insts;
    EXCEPTION_CODE         pipeline_error_status;
    logic [4:0]            pipeline_commit_wr_idx;
    logic [`XLEN-1:0]      pipeline_commit_wr_data;
    logic                   pipeline_commit_wr_en;
    logic [`XLEN-1:0]      pipeline_commit_NPC;
    logic [`XLEN-1:0]      if_NPC_dbg;
    logic [31:0]           if_inst_dbg;
    logic                   if_valid_dbg;
    logic [`XLEN-1:0]      ex_mem_NPC_dbg;
    logic [31:0]           ex_mem_inst_dbg;
    logic                   ex_mem_valid_dbg;
    logic [`XLEN-1:0]      mem_wb_NPC_dbg;
    logic [31:0]           mem_wb_inst_dbg;
    logic                   mem_wb_valid_dbg;
    MAP_PACKET [31:0]      m_table_dbg;
    logic [`NUM_FU:0]      dones_dbg;
    logic [`NUM_FU:0]      ack_dbg;
    CDB_PACKET             cdb_packet_dbg;
    CDB_EX_PACKET          cdb_ex_packet_dbg;
    MAP_RS_PACKET          map_rs_packet_dbg;
    MAP_ROB_PACKET         map_rob_packet_dbg;
    EX_CDB_PACKET          ex_cdb_packet_dbg;
    DP_PACKET              dp_packet_dbg;
    logic                  dp_packet_req_dbg;
    RS_DP_PACKET           avail_vec_dbg;
    RS_EX_PACKET           rs_ex_packet_dbg;
    ROB_RS_PACKET          rob_rs_packet_dbg;
    ROB_MAP_PACKET         rob_map_packet_dbg;
    logic                  rob_dp_available_dbg;
    ROB_RT_PACKET          rob_rt_packet_dbg;
    logic                  dispatch_valid_dbg;
    logic [`XLEN-1:0]      id_ex_inst_dbg;
    RT_DP_PACKET           rt_dp_packet_dbg;
    IB_DP_PACKET           ib_dp_packet_dbg;
    IF_IB_PACKET           if_ib_packet_dbg;
    logic                  ib_full_dbg;
    logic                  ib_empty_dbg;
    logic                  squash_dbg;

    // Instantiate the Pipeline
    pipeline pipeline_0 (
        // Inputs
        .clock             (clock),
        .reset             (reset),
        .mem2proc_response (mem2proc_response),
        .mem2proc_data     (mem2proc_data),
        .mem2proc_tag      (mem2proc_tag),

        // Outputs
        .proc2mem_command (proc2mem_command),
        .proc2mem_addr    (proc2mem_addr),
        .proc2mem_data    (proc2mem_data),
        .proc2mem_size    (proc2mem_size),

        .pipeline_completed_insts (pipeline_completed_insts),
        .pipeline_error_status    (pipeline_error_status),
        .pipeline_commit_wr_data  (pipeline_commit_wr_data),
        .pipeline_commit_wr_idx   (pipeline_commit_wr_idx),
        .pipeline_commit_wr_en    (pipeline_commit_wr_en),
        .pipeline_commit_NPC      (pipeline_commit_NPC),

        .if_NPC_dbg       (if_NPC_dbg),
        .if_inst_dbg      (if_inst_dbg),
        .if_valid_dbg     (if_valid_dbg),
        .ex_mem_NPC_dbg   (ex_mem_NPC_dbg),
	.ex_mem_inst_dbg  (ex_mem_inst_dbg),
	.ex_mem_valid_dbg (ex_mem_valid_dbg),
	.mem_wb_NPC_dbg   (mem_wb_NPC_dbg),
	.mem_wb_inst_dbg  (mem_wb_inst_dbg),
	.mem_wb_valid_dbg (mem_wb_valid_dbg),
	.m_table_dbg      (m_table_dbg),
	.dones_dbg        (dones_dbg),
	.ack_dbg          (ack_dbg),
	.cdb_packet_dbg	  (cdb_packet_dbg),
	.cdb_ex_packet_dbg(cdb_ex_packet_dbg),
	.map_rs_packet_dbg(map_rs_packet_dbg),
	.map_rob_packet_dbg    (map_rob_packet_dbg),
	.ex_cdb_packet_dbg     (ex_cdb_packet_dbg),
	.dp_packet_dbg         (dp_packet_dbg),
	.dp_packet_req_dbg     (dp_packet_req_dbg),
	.avail_vec_dbg         (avail_vec_dbg),
	.rs_ex_packet_dbg      (rs_ex_packet_dbg),
	.rob_rs_packet_dbg     (rob_rs_packet_dbg),
	.rob_map_packet_dbg    (rob_map_packet_dbg),
	.rob_dp_available_dbg  (rob_dp_available_dbg),
	.rob_rt_packet_dbg     (rob_rt_packet_dbg),
	.dispatch_valid_dbg    (dispatch_valid_dbg),
	.id_ex_inst_dbg        (id_ex_inst_dbg),
	.rt_dp_packet_dbg      (rt_dp_packet_dbg),
	.ib_dp_packet_dbg      (ib_dp_packet_dbg),
	.if_ib_packet_dbg      (if_ib_packet_dbg),
	.ib_full_dbg           (ib_full_dbg),
	.ib_empty_dbg          (ib_empty_dbg),
	.squash_dbg            (squash_dbg)
	
    );

    // Instantiate the Data Memory
    mem memory (
        // Inputs
        .clk              (clock),
        .proc2mem_command (proc2mem_command),
        .proc2mem_addr    (proc2mem_addr),
        .proc2mem_data    (proc2mem_data),
`ifndef CACHE_MODE
        .proc2mem_size    (proc2mem_size),
`endif

        // Outputs
        .mem2proc_response (mem2proc_response),
        .mem2proc_data     (mem2proc_data),
        .mem2proc_tag      (mem2proc_tag)																																																																																																																																																																																														
    );


    // Generate System Clock
    always begin
    #(`CLOCK_PERIOD/2.0);
        clock = ~clock;
    end


    // Count the number of posedges and number of instructions completed
    // till simulation ends
    always @(posedge clock) begin
        if (reset) begin
            clock_count <= 0;
            instr_count <= 0;
        end else begin
            clock_count <= (clock_count + 1);
            instr_count <= (instr_count + pipeline_completed_insts);
        end
    end


    initial begin
        clock = 0;
        reset = 0;

        // Call to initialize visual debugger
        // *Note that after this, all stdout output goes to visual debugger*
        // each argument is number of registers/signals for the group
       initcurses(
            5,  // IF
            23,  // IB
            22, // DP
            40, // RS
            48,  // MT 
            48,  // ROB
            22,  // EX
            2,  // CDB
            3,  // GLOBAL
            0   // Miscellaneous
        );

        // Pulse the reset signal
        reset = 1'b1;
        @(posedge clock);
        @(posedge clock);

        // set paramterized strings, see comment at start of module
        if ($value$plusargs("MEMORY=%s", program_memory_file)) begin
            $display("Loading memory file: %s", program_memory_file);
        end else begin
            $display("Loading default memory file: program.mem");
            program_memory_file = "program.mem";
        end

        // Read program contents into memory array
        $readmemh(program_memory_file, memory.unified_memory);
        @(posedge clock);
        @(posedge clock);
        #1;
        // This reset is at an odd time to avoid the pos & neg clock edges
        reset = 1'b0;
    end


    always @(negedge clock) begin
        if (!reset) begin
            #2;

            // deal with any halting conditions
            if (pipeline_error_status!=NO_ERROR) begin
                #100
                $display("\nDONE\n");
                waitforresponse();
                flushpipe();
                $finish;
            end
        end
    end 


    // This block is where we dump all of the signals that we care about to
    // the visual debugger.  Notice this happens at *every* clock edge.
    always @(clock) begin
        #2;

        // Dump clock and time onto stdout
        $display("c%h%7.0d",clock,clock_count);
        $display("t%8.0f",$time);
        $display("z%h",reset);

        // Dump register file contents
        $write("a");
        for(int i = 0; i < 32; i=i+1) begin
            $write("%h", pipeline_0.u_stage_dp.regfile.registers[i]);
        end
        $display("");

        // Dump instructions and their validity for each stage
        $write("p");
        $write("%h%h ",
               if_inst_dbg,      if_valid_dbg,
               );
        $display("");

        // Dump interesting register/signal contents onto stdout
        // format is "<reg group prefix><name> <width in hex chars>:<data>"
        // Current register groups (and prefixes) are:
        // f: IF   d: ID   e: EX   m: MEM    w: WB  v: misc. reg
        // g: IF/ID   h: ID/EX  i: EX/MEM  j: MEM/WB

        // IF signals (5) - prefix 'f'
        $display("finst 8:%h",        pipeline_0.if_ib_packet.inst);
	$display("fPC 8:%h",          pipeline_0.if_ib_packet.PC);
	$display("fNPC 8:%h",         pipeline_0.if_ib_packet.NPC);
        $display("fvalid 1:%h",       pipeline_0.if_ib_packet.valid);
	$display("fImem_addr 8:%h",   pipeline_0.proc2Imem_addr);

        // IB signals (4) - prefix 'g'
        
        $display("ginst 8:%h",        pipeline_0.ib_dp_packet.inst);
        $display("gPC 8:%h",          pipeline_0.ib_dp_packet.PC);
	$display("gNPC 8:%h",         pipeline_0.ib_dp_packet.NPC);
        $display("gvalid 1:%h",       pipeline_0.ib_dp_packet.valid);
	$display("gib_full 1:%h",     pipeline_0.ib_full);
        $display("gib_empty 1:%h",    pipeline_0.ib_empty);
	$display("gIB_BUFFER");
	$display("ge0 8:%h",      pipeline_0.u_insn_buffer.buffer[0].PC);
	$display("ge1 8:%h",      pipeline_0.u_insn_buffer.buffer[1].PC);
	$display("ge2 8:%h",      pipeline_0.u_insn_buffer.buffer[2].PC);
	$display("ge3 8:%h",      pipeline_0.u_insn_buffer.buffer[3].PC);
	$display("ge4 8:%h",      pipeline_0.u_insn_buffer.buffer[4].PC);
	$display("ge5 8:%h",      pipeline_0.u_insn_buffer.buffer[5].PC);
	$display("ge6 8:%h",      pipeline_0.u_insn_buffer.buffer[6].PC);
	$display("ge7 8:%h",      pipeline_0.u_insn_buffer.buffer[7].PC);
	$display("ge8 8:%h",      pipeline_0.u_insn_buffer.buffer[8].PC);
	$display("ge9 8:%h",      pipeline_0.u_insn_buffer.buffer[9].PC);
	$display("ge10 8:%h",      pipeline_0.u_insn_buffer.buffer[10].PC);
	$display("ge11 8:%h",      pipeline_0.u_insn_buffer.buffer[11].PC);
	$display("ge12 8:%h",      pipeline_0.u_insn_buffer.buffer[12].PC);
	$display("ge13 8:%h",      pipeline_0.u_insn_buffer.buffer[13].PC);
	$display("ge14 8:%h",      pipeline_0.u_insn_buffer.buffer[14].PC);
	$display("ge15 8:%h",      pipeline_0.u_insn_buffer.buffer[15].PC);



        // DP signals (13) - prefix 'd'
        $display("dfu_sel 1:%h",     		pipeline_0.dp_packet.fu_sel);
        $display("dinst 8:%h",       		pipeline_0.dp_packet.inst);
        $display("dPC 8:%h",         		pipeline_0.dp_packet.PC);
        $display("dNPC 8:%h",         		pipeline_0.dp_packet.NPC);
        $display("drs1_value 8:%h",  		pipeline_0.dp_packet.rs1_value);
        $display("drs2_value 8:%h",  		pipeline_0.dp_packet.rs2_value);
        $display("drs1_idx 2:%h",    		pipeline_0.dp_packet.rs1_idx);
        $display("drs1_idx 2:%h",    		pipeline_0.dp_packet.rs2_idx);
        $display("drs1_valid 1:%h",  		pipeline_0.dp_packet.rs1_valid); 
        $display("drs2_valid 1:%h",  		pipeline_0.dp_packet.rs2_valid);
        $display("dopa_select 1:%h", 		pipeline_0.dp_packet.opa_select);
        $display("dopb_select 1:%h", 		pipeline_0.dp_packet.opb_select);
        $display("ddest_reg_idx 2:%h",       	pipeline_0.dp_packet.dest_reg_idx);
	$display("dhas_dest 1:%h",     	pipeline_0.dp_packet.has_dest);
        $display("dalu_func 2:%h",       	pipeline_0.dp_packet.alu_func);
        $display("drd_mem 1:%h",         	pipeline_0.dp_packet.rd_mem);
        $display("dwr_mem 1:%h",         	pipeline_0.dp_packet.wr_mem);
        $display("dcond_branch 1:%h",  	pipeline_0.dp_packet.cond_branch);
        $display("duncond_branch 1:%h",  	pipeline_0.dp_packet.uncond_branch);
        $display("dhalt 1:%h",    		pipeline_0.dp_packet.halt);
        $display("dillegal 1:%h",    		pipeline_0.dp_packet.illegal);
        $display("dcsr_op 1:%h",  		pipeline_0.dp_packet.csr_op);

        // RS signals (17) - prefix 'h'
	$display("he2_fu 1:%h",      	pipeline_0.u_rs.entry[2].fu);
        $display("he2_busy 1:%h",      	pipeline_0.u_rs.entry[2].busy);
	$display("he2_r 4:%b",      	pipeline_0.u_rs.entry[2].r);
	$display("he2_t1 4:%b",      	pipeline_0.u_rs.entry[2].t1);
	$display("he2_t2 4:%b",      	pipeline_0.u_rs.entry[2].t2);
	$display("he2_v1 8:%h",      	pipeline_0.u_rs.entry[2].v1);
	$display("he2_v2 8:%h",      	pipeline_0.u_rs.entry[2].v2);
	$display("he2_issued 1:%h",     pipeline_0.u_rs.entry[2].issued);

	$display("he3_fu 1:%h",      	pipeline_0.u_rs.entry[3].fu);
        $display("he3_busy 1:%h",      	pipeline_0.u_rs.entry[3].busy);
	$display("he3_r 4:%b",      	pipeline_0.u_rs.entry[3].r);
	$display("he3_t1 4:%b",      	pipeline_0.u_rs.entry[3].t1);
	$display("he3_t2 4:%b",      	pipeline_0.u_rs.entry[3].t2);
	$display("he3_v1 8:%h",      	pipeline_0.u_rs.entry[3].v1);
	$display("he3_v2 8:%h",      	pipeline_0.u_rs.entry[3].v2);
	$display("he3_issued 1:%h",     pipeline_0.u_rs.entry[3].issued);

	$display("he4_fu 1:%h",      	pipeline_0.u_rs.entry[4].fu);
        $display("he4_busy 1:%h",      	pipeline_0.u_rs.entry[4].busy);
	$display("he4_r 4:%b",      	pipeline_0.u_rs.entry[4].r);
	$display("he4_t1 4:%b",      	pipeline_0.u_rs.entry[4].t1);
	$display("he4_t2 4:%b",      	pipeline_0.u_rs.entry[4].t2);
	$display("he4_v1 8:%h",      	pipeline_0.u_rs.entry[4].v1);
	$display("he4_v2 8:%h",      	pipeline_0.u_rs.entry[4].v2);
	$display("he4_issued 1:%h",     pipeline_0.u_rs.entry[4].issued);

	$display("he5_fu 1:%h",      	pipeline_0.u_rs.entry[5].fu);
        $display("he5_busy 1:%h",      	pipeline_0.u_rs.entry[5].busy);
	$display("he5_r 4:%b",      	pipeline_0.u_rs.entry[5].r);
	$display("he5_t1 4:%b",      	pipeline_0.u_rs.entry[5].t1);
	$display("he5_t2 4:%b",      	pipeline_0.u_rs.entry[5].t2);
	$display("he5_v1 8:%h",      	pipeline_0.u_rs.entry[5].v1);
	$display("he5_v2 8:%h",      	pipeline_0.u_rs.entry[5].v2);
	$display("he5_issued 1:%h",     pipeline_0.u_rs.entry[5].issued);


	$display("he6_fu 1:%h",      	pipeline_0.u_rs.entry[6].fu);
        $display("he6_busy 1:%h",      	pipeline_0.u_rs.entry[6].busy);
	$display("he6_r 4:%b",      	pipeline_0.u_rs.entry[6].r);
	$display("he6_t1 4:%b",      	pipeline_0.u_rs.entry[6].t1);
	$display("he6_t2 4:%b",      	pipeline_0.u_rs.entry[6].t2);
	$display("he6_v1 8:%h",      	pipeline_0.u_rs.entry[6].v1);
	$display("he6_v2 8:%h",       	pipeline_0.u_rs.entry[6].v2);
	$display("he6_issued 1:%h",     pipeline_0.u_rs.entry[6].issued);

        // MT signals (4) - prefix 'e'
	$display("ee0 4:%b",     pipeline_0.u_map_table.m_table[0].rob_tag);
	$display("ee0 1:%b",     pipeline_0.u_map_table.m_table[0].t_plus);
        $display("ee1 4:%b",     pipeline_0.u_map_table.m_table[1].rob_tag);
	$display("ee1 1:%b",     pipeline_0.u_map_table.m_table[1].t_plus);
	$display("ee2 4:%b",     pipeline_0.u_map_table.m_table[2].rob_tag);
	$display("ee2 1:%b",     pipeline_0.u_map_table.m_table[2].t_plus);
	$display("ee3 4:%b",     pipeline_0.u_map_table.m_table[3].rob_tag);
	$display("ee3 1:%b",     pipeline_0.u_map_table.m_table[3].t_plus);
	$display("ee4 4:%b",     pipeline_0.u_map_table.m_table[4].rob_tag);
	$display("ee4 1:%b",     pipeline_0.u_map_table.m_table[4].t_plus);
	$display("ee5 4:%b",     pipeline_0.u_map_table.m_table[5].rob_tag);
	$display("ee5 1:%b",     pipeline_0.u_map_table.m_table[5].t_plus);
        $display("ee6 4:%b",     pipeline_0.u_map_table.m_table[6].rob_tag);
	$display("ee6 1:%b",     pipeline_0.u_map_table.m_table[6].t_plus);
	$display("ee7 4:%b",     pipeline_0.u_map_table.m_table[7].rob_tag);
	$display("ee7 1:%b",     pipeline_0.u_map_table.m_table[7].t_plus);
	$display("ee8 4:%b",     pipeline_0.u_map_table.m_table[8].rob_tag);
	$display("ee8 1:%b",     pipeline_0.u_map_table.m_table[8].t_plus);
	$display("ee9 4:%b",     pipeline_0.u_map_table.m_table[9].rob_tag);
	$display("ee9 1:%b",     pipeline_0.u_map_table.m_table[9].t_plus);
	$display("ee10 4:%b",     pipeline_0.u_map_table.m_table[10].rob_tag);
	$display("ee10 1:%b",     pipeline_0.u_map_table.m_table[10].t_plus);
        $display("ee11 4:%b",     pipeline_0.u_map_table.m_table[11].rob_tag);
	$display("ee11 1:%b",     pipeline_0.u_map_table.m_table[11].t_plus);
	$display("ee12 4:%b",     pipeline_0.u_map_table.m_table[12].rob_tag);
	$display("ee12 1:%b",     pipeline_0.u_map_table.m_table[12].t_plus);
	$display("ee13 4:%b",     pipeline_0.u_map_table.m_table[13].rob_tag);
	$display("ee13 1:%b",     pipeline_0.u_map_table.m_table[13].t_plus);
	$display("ee14 4:%b",     pipeline_0.u_map_table.m_table[14].rob_tag);
	$display("ee14 1:%b",     pipeline_0.u_map_table.m_table[14].t_plus);	
	$display("ee15 4:%b",     pipeline_0.u_map_table.m_table[15].rob_tag);
	$display("ee15 1:%b",     pipeline_0.u_map_table.m_table[15].t_plus);
        $display("ee16 4:%b",     pipeline_0.u_map_table.m_table[16].rob_tag);
	$display("ee16 1:%b",     pipeline_0.u_map_table.m_table[16].t_plus);
	$display("ee17 4:%b",     pipeline_0.u_map_table.m_table[17].rob_tag);
	$display("ee17 1:%b",     pipeline_0.u_map_table.m_table[17].t_plus);
	$display("ee18 4:%b",     pipeline_0.u_map_table.m_table[18].rob_tag);
	$display("ee18 1:%b",     pipeline_0.u_map_table.m_table[18].t_plus);
	$display("ee19 4:%b",     pipeline_0.u_map_table.m_table[19].rob_tag);
	$display("ee19 1:%b",     pipeline_0.u_map_table.m_table[19].t_plus);
	$display("ee20 4:%b",     pipeline_0.u_map_table.m_table[20].rob_tag);
	$display("ee20 1:%b",     pipeline_0.u_map_table.m_table[20].t_plus);
        $display("ee21 4:%b",     pipeline_0.u_map_table.m_table[21].rob_tag);
	$display("ee21 1:%b",     pipeline_0.u_map_table.m_table[21].t_plus);
	$display("ee22 4:%b",     pipeline_0.u_map_table.m_table[22].rob_tag);
	$display("ee22 1:%b",     pipeline_0.u_map_table.m_table[22].t_plus);
	$display("ee23 4:%b",     pipeline_0.u_map_table.m_table[23].rob_tag);
	$display("ee23 1:%b",     pipeline_0.u_map_table.m_table[23].t_plus);
	
        
        // ROB signals (14) - prefix 'i'
	$display("ie24 4:%b",     pipeline_0.u_map_table.m_table[24].rob_tag);
	$display("ie24 1:%b",     pipeline_0.u_map_table.m_table[24].t_plus);
	$display("ie25 4:%b",     pipeline_0.u_map_table.m_table[25].rob_tag);
	$display("ie25 1:%b",     pipeline_0.u_map_table.m_table[25].t_plus);
	$display("ie26 4:%b",     pipeline_0.u_map_table.m_table[26].rob_tag);
	$display("ie26 1:%b",     pipeline_0.u_map_table.m_table[26].t_plus);
	$display("ie27 4:%b",     pipeline_0.u_map_table.m_table[27].rob_tag);
	$display("ie27 1:%b",     pipeline_0.u_map_table.m_table[27].t_plus);
	$display("ie28 4:%b",     pipeline_0.u_map_table.m_table[28].rob_tag);
	$display("ie28 1:%b",     pipeline_0.u_map_table.m_table[28].t_plus);
	$display("ie29 4:%b",     pipeline_0.u_map_table.m_table[29].rob_tag);
	$display("ie29 1:%b",     pipeline_0.u_map_table.m_table[29].t_plus);
	$display("ie30 4:%b",     pipeline_0.u_map_table.m_table[30].rob_tag);
	$display("ie30 1:%b",     pipeline_0.u_map_table.m_table[30].t_plus);
	$display("ie31 4:%b",     pipeline_0.u_map_table.m_table[31].rob_tag);
	$display("ie31 1:%b",     pipeline_0.u_map_table.m_table[31].t_plus);

	$display("ie1_r 5:%b",      pipeline_0.u_rob.rob_memory[1].r);
	$display("ie1_V 8:%h",      pipeline_0.u_rob.rob_memory[1].V);
	$display("ie1_rob_tag 4:%b",pipeline_0.u_rob.rob_memory[1].rob_tag);
	$display("ie1_done 1:%b",      pipeline_0.u_rob.rob_memory[1].complete);
	$display("ie2_r 5:%b",      pipeline_0.u_rob.rob_memory[2].r);
	$display("ie2_V 8:%h",      pipeline_0.u_rob.rob_memory[2].V);
	$display("ie2_rob_tag 4:%b",pipeline_0.u_rob.rob_memory[2].rob_tag);
	$display("ie2_done 1:%b",      pipeline_0.u_rob.rob_memory[2].complete);
	$display("ie3_r 5:%b",      pipeline_0.u_rob.rob_memory[3].r);
	$display("ie3_V 8:%h",      pipeline_0.u_rob.rob_memory[3].V);
	$display("ie3_rob_tag 4:%b",pipeline_0.u_rob.rob_memory[3].rob_tag);
	$display("ie3_done 1:%b",      pipeline_0.u_rob.rob_memory[3].complete);
	$display("ie4_r 5:%b",      pipeline_0.u_rob.rob_memory[4].r);
	$display("ie4_V 8:%h",      pipeline_0.u_rob.rob_memory[4].V);
	$display("ie4_rob_tag 4:%b",pipeline_0.u_rob.rob_memory[4].rob_tag);
	$display("ie4_done 1:%b",      pipeline_0.u_rob.rob_memory[4].complete);
	$display("ie5_r 5:%b",      pipeline_0.u_rob.rob_memory[5].r);
	$display("ie5_V 8:%h",      pipeline_0.u_rob.rob_memory[5].V);
	$display("ie5_rob_tag 4:%b",pipeline_0.u_rob.rob_memory[5].rob_tag);
	$display("ie5_done 1:%b",      pipeline_0.u_rob.rob_memory[5].complete);
	$display("ie6_r 5:%b",      pipeline_0.u_rob.rob_memory[6].r);
	$display("ie6_V 8:%h",      pipeline_0.u_rob.rob_memory[6].V);
	$display("ie6_rob_tag 4:%b",pipeline_0.u_rob.rob_memory[6].rob_tag);
	$display("ie6_done 1:%b",      pipeline_0.u_rob.rob_memory[6].complete);
	$display("ie7_r 5:%b",      pipeline_0.u_rob.rob_memory[7].r);
	$display("ie7_V 8:%h",      pipeline_0.u_rob.rob_memory[7].V);
	$display("ie7_rob_tag 4:%b",pipeline_0.u_rob.rob_memory[7].rob_tag);
	$display("ie7_done 1:%b",      pipeline_0.u_rob.rob_memory[7].complete);
	$display("ie8_r 5:%b",      pipeline_0.u_rob.rob_memory[8].r);
	$display("ie8_V 8:%h",      pipeline_0.u_rob.rob_memory[8].V);
	$display("ie8_rob_tag 4:%b",pipeline_0.u_rob.rob_memory[8].rob_tag);
	$display("ie8_done 1:%b",      pipeline_0.u_rob.rob_memory[8].complete);

        // EX signals (5) - prefix 'm'
	$display("me0_r 5:%b",      pipeline_0.u_rob.rob_memory[0].r);
	$display("me0_V 8:%h",      pipeline_0.u_rob.rob_memory[0].V);
	$display("me0_rob_tag 4:%b",pipeline_0.u_rob.rob_memory[0].rob_tag);
	$display("me0_done 1:%b",      pipeline_0.u_rob.rob_memory[0].complete);
        $display("malu1_done 1:%h",   	pipeline_0.u_ex.fu_1.fu_out_packet.done);
        $display("malu1_v 8:%h",  	pipeline_0.u_ex.fu_1.fu_out_packet.v);
	$display("malu1_robtag 4:%b",  	pipeline_0.u_ex.fu_1.fu_out_packet.rob_tag);
	$display("malu2_done 1:%h",   	pipeline_0.u_ex.fu_2.fu_out_packet.done);
        $display("malu2_v 8:%h",  	pipeline_0.u_ex.fu_2.fu_out_packet.v);
	$display("malu2_robtag 4:%b",  	pipeline_0.u_ex.fu_2.fu_out_packet.rob_tag);
	$display("mload_done 1:%h",   	pipeline_0.u_ex.fu_3.fu_out_packet.done);
        $display("mload_v 8:%h",  	pipeline_0.u_ex.fu_3.fu_out_packet.v);
	$display("mload_robtag 4:%b",  	pipeline_0.u_ex.fu_3.fu_out_packet.rob_tag);
	$display("mstore_done 1:%h",   	pipeline_0.u_ex.fu_4.fu_out_packet.done);
        $display("mstore_v 8:%h",  	pipeline_0.u_ex.fu_4.fu_out_packet.v);
	$display("mstore_robtag 4:%b",  pipeline_0.u_ex.fu_4.fu_out_packet.rob_tag);
	$display("mmult1_done 1:%h",   	pipeline_0.u_ex.fu_5.fu_out_packet.done);
        $display("mmult1_v 8:%h",  	pipeline_0.u_ex.fu_5.fu_out_packet.v);
	$display("mmult1_robtag 4:%b",  pipeline_0.u_ex.fu_5.fu_out_packet.rob_tag);
	$display("mmult2_done 1:%h",   	pipeline_0.u_ex.fu_6.fu_out_packet.done);
        $display("mmult2_v 8:%h",  	pipeline_0.u_ex.fu_6.fu_out_packet.v);
	$display("mmult2_robtag 4:%b",  pipeline_0.u_ex.fu_6.fu_out_packet.rob_tag);
	
      

        // CDB signals (9) - prefix 'j'
        $display("jrob_tag 4:%b",      pipeline_0.cdb_packet.rob_tag);
        $display("jv 8:%h",            pipeline_0.cdb_packet.v);
        

        // GLOBAL signals (3) - prefix 'w'
        $display("wdispatch_valid 1:%h",     pipeline_0.dispatch_valid);
        $display("wsquash 1:%h",      pipeline_0.squash);
        $display("wreset 1:%h",       pipeline_0.reset); 

        // Misc signals(2) - prefix 'v'
        /*$display("vcompleted 1:%h",   pipeline_completed_insts);
        $display("vpipe_err 1:%h",    pipeline_error_status); */

        // must come last
        $display("break");

        // This is a blocking call to allow the debugger to control when we
        // advance the simulation
        waitforresponse();
    end

endmodule // module testbench
